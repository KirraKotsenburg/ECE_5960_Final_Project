/*********************
El Gamal Circuit (Toplevel)
contains encrypt and decrypt
*********************/
module ElGamal(

);

endmodule