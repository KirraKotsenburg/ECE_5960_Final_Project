module encrypt(
		input [3:0] e1x,
		input [3:0] e1y,
		input [3:0] e1z,
		input [3:0] e2x,
		input [3:0] e2y,
		input [3:0] e2z,
		input [3:0] Epx,
		input [3:0] Epy,
		input [3:0] EpZ,
		output [3:0] C1x,
		output [3:0] C1y,
		output [3:0] C1z,
		output [3:0] C2x,
		output [3:0] C2y,
		output [3:0] C2z

);

endmodule
