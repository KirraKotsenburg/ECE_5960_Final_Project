
module pointADD(

);


endmodule