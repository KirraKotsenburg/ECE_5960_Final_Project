module decrypt(

);


endmodule