/*********************
El Gamal Circuit (Toplevel)
contains encrypt and decrypt
Key genration module inside as well
*********************/
module ElGamal(

);

endmodule