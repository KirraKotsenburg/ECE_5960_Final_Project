
module pointDouble(

);


endmodule