module keygen(

);


endmodule
