`include "control_if.vh"    

module control (
  input logic nRST,
  control_if.co coif
);
  
  always_comb begin 
    
  end
endmodule