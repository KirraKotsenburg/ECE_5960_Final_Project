module 4b_MMult(
    input [3:0]A,
    input [3:0] B,
    output reg[3:0] Z
    );

// Temporary reg
reg [6:0] S;

always@(*) begin
    
    


end

endmodule 