`timescale 1ps/1ps

module pointAdd (
  input logic[3:0] X0, Y0, Z0, X1, Y1, Z1,
  output logic[3:0] X2, Y2, Z2
);
  logic[3:0] A0, A1, B0, B1, C, D, E, F, G, H, I, J;

  MMult

  always_comb begin
    A0 = 
  end


endmodule