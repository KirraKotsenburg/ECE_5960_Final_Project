/*********************
Key Generation for El Gamal
Selection for d, e1, Ep
e2 needs to be calculated
*********************/
module keygen(

);


endmodule
