module encrypt(

);

endmodule
